// alu.v
// ECE 154A, Fall 2019
// Authors: Daniel Kluzner, Benji

// A 32-bit arithmetic logic unit (ALU)
// as seen in 5.2.4 of "Harris & Harris"

module alu(
       input [31:0] a,
       input [31:0] b,
       input [2:0] f,
       output [31:0] y,
       output zero
);

// CODE

endmodule
