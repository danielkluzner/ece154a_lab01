// testbench.v
// ECE 154A, Fall 2019
// Authors: Daniel Kluzner, Benji

// A testbench for the "alu" module

module alu_tb();

// CODE

endmodule

